`timescale 1ns / 1ps

module tb_CPU( );

    integer i = 1;
    integer j = 0;
    
    
    reg clk, rstn, cnt_start;
    reg [7:0] memory_8 [0:511];
    
    CPU_top uut(clk,rstn);
    
    always@(posedge clk)
        if(cnt_start) j <= j + 1;
    
    initial begin 
        memory_8[0:79] = 
        {
            8'b00000000, 8'b00100000, 8'b10000000, 8'b10010011, //     addi x1, x1, #2
            8'b00000000, 8'b00100011, 8'b00000011, 8'b01111111, //     illegal opcode
            8'b00010000, 8'b00010001, 8'b10000001, 8'b10010011, //     addi x3, x3, #101
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, //
            8'b00010000, 8'b00010010, 8'b00000010, 8'b00010011, //     addi x4, x4, #101
            8'b00111110, 8'b10000010, 8'b10100101, 8'b00000011, //     lw x10, [x5, #d'1000] (load/store access fault)
            8'b00010000, 8'b00010001, 8'b10000001, 8'b10010011, //     addi x3, x3, #101
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, //
            8'b00010000, 8'b00010010, 8'b00000010, 8'b00010011, //     addi x4, x4, #101
            8'b00111110, 8'b10000000, 8'b00000000, 8'b01101111, //     jal xzr, #d'1000 (instruction access fault)
            8'b00010000, 8'b00010001, 8'b10000001, 8'b10010011, //     addi x3, x3, #101
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, //
            8'b00010000, 8'b00010010, 8'b00000010, 8'b00010011, //     addi x4, x4, #101
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000,
            8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000  //       NOP


            };
            
        for(i = 80; i<472; i = i + 1) begin
            memory_8[i] = 8'b0;
        end
        
        //exception handler
        memory_8[472:511] =    
        {   //load/store access fault
            8'b00000000, 8'b00010000, 8'b10000011, 8'b10010011, //     addi x7, x1, #1
            8'b00110000, 8'b00100000, 8'b00000000, 8'b01110011, //     mret
            //illegal instruction
            8'b00000000, 8'b00100000, 8'b10000011, 8'b10010011, //     addi x7, x1, #2
            8'b00110000, 8'b00100000, 8'b00000000, 8'b01110011, //     mret
            //instruction access fault
            8'b00000000, 8'b00110000, 8'b10000011, 8'b10010011, //     addi x7, x1, #3
            8'b00110000, 8'b00100000, 8'b00000000, 8'b01110011, //     mret
            //--------------------------------------------------------------------------------------
            8'b00000000, 8'b00100000, 8'b10000011, 8'b10010011, //     addi x7, x1, #2
            8'b00110000, 8'b00100000, 8'b00000000, 8'b01110011, //     mret
            8'b00000000, 8'b00100000, 8'b10000011, 8'b10010011, //     addi x7, x1, #2
            8'b00110000, 8'b00100000, 8'b00000000, 8'b01110011 //     mret
            };
    end
    
    initial begin
        for(i = 0; i<128; i = i+1)begin
            uut.instruction_cache_mem.inst_mem_L1[i] = 
                {memory_8[4*i],memory_8[4*i+1],memory_8[4*i+2],memory_8[4*i+3]};
        end
    end
    
    initial begin 
        clk = 0;
        forever #5 clk = ~clk;
    end
    
    initial begin
        cnt_start = 0;
        rstn = 0;
        
        #25
        rstn = 1;
        
        #10
        cnt_start = 1;
    end
    
    initial #2000 $finish;

endmodule
